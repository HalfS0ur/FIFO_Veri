//Second